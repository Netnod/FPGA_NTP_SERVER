module ntps_top_axi_ethernetlite_0_0 (
    input wire         s_axi_aclk,
    input wire         s_axi_aresetn,
    output wire        ip2intc_irpt,
    input wire [12:0]  s_axi_awaddr,
    input wire         s_axi_awvalid,
    output wire        s_axi_awready,
    input wire [31:0]  s_axi_wdata,
    input wire [3:0]   s_axi_wstrb,
    input wire         s_axi_wvalid,
    output wire        s_axi_wready,
    output wire [1:0]  s_axi_bresp,
    output wire        s_axi_bvalid,
    input wire         s_axi_bready,
    input wire [12:0]  s_axi_araddr,
    input wire         s_axi_arvalid,
    output wire        s_axi_arready,
    output wire [31:0] s_axi_rdata,
    output wire [1:0]  s_axi_rresp,
    output wire        s_axi_rvalid,
    input wire         s_axi_rready,
    input wire         phy_tx_clk,
    input wire         phy_rx_clk,
    input wire         phy_crs,
    input wire         phy_dv,
    input wire [3:0]   phy_rx_data,
    input wire         phy_col,
    input wire         phy_rx_er,
    output wire        phy_rst_n,
    output wire        phy_tx_en,
    output wire [3:0]  phy_tx_data,
    input wire         phy_mdio_i,
    output wire        phy_mdio_o,
    output wire        phy_mdio_t,
    output wire        phy_mdc
  );
endmodule // ntps_top_axi_ethernetlite_0_0

