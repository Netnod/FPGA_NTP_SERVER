module ntps_top_clock_control_0_0 (
  inout wire  i2c_clk,
  inout wire  i2c_data,
  output wire i2c_mux_rst_n,
  output wire si5324_rst_n,
  input wire  rst,
  input wire  clk50
 );
endmodule // ntps_top_clock_control_0_0

  

