module VCC (output wire P);
  assign P = 1'b1;
endmodule // VCC

module GND (output wire G);
  assign G = 1'b0;
endmodule // GND

module ntps_top_xlconstant_0_0 (output wire [0:0] dout);
  assign dout = 1'b0;
endmodule // ntps_top_xlconstant_0_0

module ntps_top_xlconstant_1_0 (output wire [3:0] dout);
  assign dout = 4'b0;
endmodule // ntps_top_xlconstant_0_0

module ntps_top_xlconstant_0_1 (output wire [0:0] dout);
  assign dout = 1'b0;
endmodule // ntps_top_xlconstant_0_0

