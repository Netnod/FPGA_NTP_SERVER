module ntps_top_util_ds_buf_0_0 (
    input wire  IBUF_DS_P,
    input wire  IBUF_DS_N,
    output wire IBUF_OUT,
    output wire IBUF_DS_ODIV2
  );
endmodule // ntps_top_util_ds_buf_0_0


